magic
tech sample_6m
timestamp 1598177544
<< nwell >>
rect -93 -33 -60 -4
rect 0 -14 23 44
rect 56 -32 89 -3
<< ntransistor >>
rect -52 -19 -48 -17
rect 44 -18 48 -16
rect 7 -29 12 -27
rect 7 -50 12 -48
<< ptransistor >>
rect 5 18 14 20
rect 5 -2 14 0
rect -76 -19 -66 -17
rect 62 -18 72 -16
<< ndiffusion >>
rect -52 -17 -48 -14
rect 44 -16 48 -13
rect -52 -22 -48 -19
rect 7 -21 12 -20
rect 44 -21 48 -18
rect 7 -27 12 -26
rect 7 -30 12 -29
rect 7 -36 12 -35
rect 7 -42 12 -41
rect 7 -48 12 -47
rect 7 -52 12 -50
<< pdiffusion >>
rect 5 26 14 27
rect 5 21 7 26
rect 12 21 14 26
rect 5 20 14 21
rect 5 17 14 18
rect 5 12 7 17
rect 12 12 14 17
rect 5 11 14 12
rect 5 6 14 7
rect 5 1 7 6
rect 12 1 14 6
rect 5 0 14 1
rect 5 -3 14 -2
rect 5 -8 7 -3
rect 12 -8 14 -3
rect 5 -9 14 -8
rect -76 -14 -71 -9
rect 67 -13 72 -8
rect -76 -17 -66 -14
rect 62 -16 72 -13
rect -76 -22 -66 -19
rect -71 -27 -66 -22
rect 62 -21 72 -18
rect 62 -26 67 -21
<< ndcontact >>
rect -53 -14 -48 -9
rect 44 -13 49 -8
rect -52 -27 -47 -22
rect 7 -26 12 -21
rect 43 -26 48 -21
rect 7 -35 12 -30
rect 7 -47 12 -42
rect 7 -57 12 -52
<< pdcontact >>
rect 7 21 12 26
rect 7 12 12 17
rect 7 1 12 6
rect 7 -8 12 -3
rect -71 -14 -66 -9
rect 62 -13 67 -8
rect -76 -27 -71 -22
rect 67 -26 72 -21
<< psubstratepcontact >>
rect -37 -14 -32 -9
rect 28 -13 33 -8
rect -37 -27 -32 -22
rect 28 -26 33 -21
rect 7 -72 12 -67
rect 17 -72 22 -67
<< nsubstratencontact >>
rect 7 37 12 42
rect 16 37 21 42
rect -91 -15 -86 -10
rect 82 -14 87 -9
rect -91 -27 -86 -22
rect 82 -26 87 -21
<< polysilicon >>
rect -2 18 5 20
rect 14 18 17 20
rect 2 -2 5 0
rect 14 -2 28 0
rect -79 -19 -76 -17
rect -66 -19 -52 -17
rect -48 -19 -45 -17
rect 41 -18 44 -16
rect 48 -18 62 -16
rect 72 -18 75 -16
rect 51 -27 53 -18
rect 4 -29 7 -27
rect 12 -29 53 -27
rect 3 -50 7 -48
rect 12 -50 15 -48
<< polycontact >>
rect -7 16 -2 21
rect 28 -4 33 1
rect -2 -51 3 -46
<< metal1 >>
rect 12 37 16 42
rect 21 37 22 42
rect 7 26 12 37
rect -59 16 -7 21
rect -59 -9 -54 16
rect -66 -14 -53 -9
rect -91 -22 -86 -15
rect -37 -22 -32 -14
rect -86 -27 -76 -22
rect -47 -27 -37 -22
rect -19 -46 -14 16
rect 7 6 12 12
rect 33 -4 55 1
rect 50 -8 55 -4
rect 7 -15 12 -8
rect 49 -13 62 -8
rect 7 -19 13 -15
rect 7 -21 12 -19
rect 28 -21 33 -13
rect 82 -21 87 -14
rect 33 -26 43 -21
rect 72 -26 82 -21
rect 7 -42 12 -35
rect -19 -51 -2 -46
rect 7 -52 12 -51
rect 7 -67 12 -57
rect 12 -72 17 -67
<< labels >>
rlabel metal1 13 -19 13 -15 1 out
rlabel polysilicon 52 -27 52 -27 1 en
rlabel metal1 14 -69 14 -69 1 gnd
rlabel metal1 13 40 13 40 5 vdd
rlabel polysilicon -57 -18 -57 -18 1 in
rlabel metal1 -89 -18 -89 -18 3 vdd
rlabel metal1 -34 -18 -34 -18 1 gnd
rlabel metal1 31 -17 31 -17 1 gnd
rlabel metal1 85 -17 85 -17 7 vdd
<< end >>
