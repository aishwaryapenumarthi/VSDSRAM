magic
tech scmos
timestamp 1598281576
<< nwell >>
rect -9 -24 15 2
rect 23 -24 43 22
rect 50 -9 74 17
<< ntransistor >>
rect 61 -19 63 -15
rect 2 -38 4 -34
rect 31 -37 35 -35
rect 31 -53 35 -51
<< ptransistor >>
rect 29 4 37 6
rect 2 -17 4 -9
rect 61 -2 63 6
rect 29 -13 37 -11
<< ndiffusion >>
rect 60 -19 61 -15
rect 63 -19 64 -15
rect 1 -38 2 -34
rect 4 -38 5 -34
rect 31 -35 35 -34
rect 31 -38 35 -37
rect 31 -51 35 -50
rect 31 -54 35 -53
<< pdiffusion >>
rect 29 7 31 11
rect 35 7 37 11
rect 29 6 37 7
rect 1 -13 2 -9
rect -3 -17 2 -13
rect 4 -13 9 -9
rect 4 -17 5 -13
rect 29 3 37 4
rect 29 -1 31 3
rect 35 -1 37 3
rect 56 2 61 6
rect 60 -2 61 2
rect 63 2 64 6
rect 63 -2 68 2
rect 29 -10 31 -6
rect 35 -10 37 -6
rect 29 -11 37 -10
rect 29 -14 37 -13
rect 29 -18 31 -14
rect 35 -18 37 -14
<< ndcontact >>
rect 56 -19 60 -15
rect 64 -19 68 -15
rect -3 -38 1 -34
rect 5 -38 9 -34
rect 31 -34 35 -30
rect 31 -42 35 -38
rect 31 -50 35 -46
rect 31 -58 35 -54
<< pdcontact >>
rect 31 7 35 11
rect -3 -13 1 -9
rect 5 -17 9 -13
rect 31 -1 35 3
rect 56 -2 60 2
rect 64 2 68 6
rect 31 -10 35 -6
rect 31 -18 35 -14
<< psubstratepcontact >>
rect 56 -29 60 -25
rect 64 -29 68 -25
rect -3 -48 1 -44
rect 5 -48 9 -44
rect 31 -66 35 -62
rect 39 -66 43 -62
<< nsubstratencontact >>
rect 26 15 30 19
rect 36 15 40 19
rect 56 10 60 14
rect 64 10 68 14
rect -3 -5 1 -1
rect 5 -5 9 -1
<< polysilicon >>
rect 61 6 63 8
rect 19 4 29 6
rect 37 4 39 6
rect 2 -9 4 -7
rect 2 -34 4 -17
rect 19 -27 21 4
rect 27 -13 29 -11
rect 37 -13 45 -11
rect 61 -11 63 -2
rect 61 -13 72 -11
rect 61 -15 63 -13
rect 61 -21 63 -19
rect 2 -40 4 -38
rect 19 -51 21 -32
rect 70 -35 72 -13
rect 29 -37 31 -35
rect 35 -37 72 -35
rect 19 -53 31 -51
rect 35 -53 37 -51
<< polycontact >>
rect 45 -14 50 -10
rect 17 -32 21 -27
<< metal1 >>
rect 30 15 36 19
rect 31 11 35 15
rect 60 10 64 14
rect 64 6 68 10
rect 1 -5 5 -1
rect -3 -9 1 -5
rect 31 -6 35 -1
rect 56 -10 60 -2
rect 50 -14 60 -10
rect 5 -27 9 -17
rect 31 -25 35 -18
rect 56 -15 60 -14
rect 64 -25 68 -19
rect 5 -32 17 -27
rect 31 -29 36 -25
rect 60 -29 64 -25
rect 31 -30 35 -29
rect 5 -34 9 -32
rect -3 -44 1 -38
rect 1 -48 5 -44
rect 31 -46 35 -42
rect 31 -62 35 -58
rect 35 -66 39 -62
<< labels >>
rlabel polysilicon 3 -30 3 -30 1 in
rlabel metal1 3 -46 3 -46 1 gnd
rlabel metal1 37 -64 37 -64 1 gnd
rlabel metal1 33 17 33 17 5 vdd
rlabel metal1 3 -3 3 -3 1 vdd
rlabel metal1 62 12 62 12 1 vdd
rlabel metal1 62 -28 62 -28 1 gnd
rlabel metal1 36 -29 36 -25 1 out
rlabel polysilicon 64 -12 64 -12 1 en
rlabel metal1 8 -29 8 -29 1 in_bar
rlabel metal1 58 -11 58 -11 1 en_bar
<< end >>
