magic
tech scmos
timestamp 1599060627
<< nwell >>
rect 1 -24 82 22
<< ntransistor >>
rect 12 -39 14 -35
rect 31 -40 35 -38
rect 51 -42 53 -38
rect 69 -40 73 -38
rect 31 -56 35 -54
rect 69 -56 73 -54
<< ptransistor >>
rect 29 4 37 6
rect 67 4 75 6
rect 12 -17 14 -9
rect 29 -12 37 -10
rect 51 -17 53 -9
rect 67 -12 75 -10
<< ndiffusion >>
rect 11 -39 12 -35
rect 14 -39 15 -35
rect 31 -38 35 -37
rect 31 -41 35 -40
rect 50 -42 51 -38
rect 53 -42 54 -38
rect 69 -38 73 -37
rect 69 -41 73 -40
rect 31 -54 35 -53
rect 69 -54 73 -53
rect 31 -57 35 -56
rect 69 -57 73 -56
<< pdiffusion >>
rect 29 7 31 11
rect 35 7 37 11
rect 29 6 37 7
rect 67 7 69 11
rect 73 7 75 11
rect 67 6 75 7
rect 29 3 37 4
rect 29 -1 31 3
rect 35 -1 37 3
rect 67 3 75 4
rect 67 -1 69 3
rect 73 -1 75 3
rect 29 -9 31 -5
rect 35 -9 37 -5
rect 67 -9 69 -5
rect 73 -9 75 -5
rect 11 -13 12 -9
rect 7 -17 12 -13
rect 14 -13 19 -9
rect 29 -10 37 -9
rect 14 -17 15 -13
rect 29 -13 37 -12
rect 46 -13 51 -9
rect 29 -17 31 -13
rect 35 -17 37 -13
rect 50 -17 51 -13
rect 53 -13 54 -9
rect 67 -10 75 -9
rect 67 -13 75 -12
rect 53 -17 58 -13
rect 67 -17 69 -13
rect 73 -17 75 -13
<< ndcontact >>
rect 7 -39 11 -35
rect 15 -39 19 -35
rect 31 -37 35 -33
rect 69 -37 73 -33
rect 31 -45 35 -41
rect 46 -42 50 -38
rect 54 -42 58 -38
rect 69 -45 73 -41
rect 31 -53 35 -49
rect 69 -53 73 -49
rect 31 -61 35 -57
rect 69 -61 73 -57
<< pdcontact >>
rect 31 7 35 11
rect 69 7 73 11
rect 31 -1 35 3
rect 69 -1 73 3
rect 31 -9 35 -5
rect 69 -9 73 -5
rect 7 -13 11 -9
rect 15 -17 19 -13
rect 31 -17 35 -13
rect 46 -17 50 -13
rect 54 -13 58 -9
rect 69 -17 73 -13
<< psubstratepcontact >>
rect 61 -61 65 -57
rect 31 -69 35 -65
<< nsubstratencontact >>
rect 31 15 35 19
rect 69 15 73 19
rect 7 -5 11 -1
rect 54 -5 58 -1
<< polysilicon >>
rect 26 4 29 6
rect 37 4 39 6
rect 65 4 67 6
rect 75 4 78 6
rect 12 -9 14 -7
rect 51 -9 53 -7
rect 27 -12 29 -10
rect 37 -12 39 -10
rect 65 -12 67 -10
rect 75 -12 77 -10
rect 12 -35 14 -17
rect 51 -26 53 -17
rect 51 -28 56 -26
rect 12 -41 14 -39
rect 29 -40 31 -38
rect 35 -40 38 -38
rect 51 -38 53 -28
rect 66 -40 69 -38
rect 73 -40 75 -38
rect 51 -44 53 -42
rect 26 -56 31 -54
rect 35 -56 37 -54
rect 67 -56 69 -54
rect 73 -56 78 -54
<< polycontact >>
rect 22 3 26 7
rect 78 3 82 7
rect 39 -13 43 -9
rect 61 -13 65 -9
rect 8 -22 12 -18
rect 38 -41 42 -37
rect 56 -29 60 -25
rect 62 -41 66 -37
rect 22 -57 26 -53
rect 78 -57 82 -53
<< metal1 >>
rect 31 11 35 15
rect 69 11 73 15
rect 11 -5 14 -1
rect 7 -9 11 -5
rect 7 -22 8 -18
rect 15 -27 19 -17
rect 22 -27 26 3
rect 31 -5 35 -1
rect 53 -5 54 -1
rect 54 -9 58 -5
rect 69 -5 73 -1
rect 15 -31 26 -27
rect 15 -35 19 -31
rect 7 -45 11 -39
rect 22 -53 26 -31
rect 31 -33 35 -17
rect 39 -25 43 -13
rect 46 -33 50 -17
rect 61 -25 65 -13
rect 60 -29 61 -25
rect 69 -33 73 -17
rect 46 -38 50 -37
rect 78 -18 82 3
rect 31 -49 35 -45
rect 54 -45 58 -42
rect 69 -49 73 -45
rect 78 -53 82 -22
rect 65 -61 69 -57
rect 31 -65 35 -61
rect 69 -65 73 -61
rect 35 -69 39 -65
<< m2contact >>
rect 35 15 39 19
rect 65 15 69 19
rect 14 -5 18 -1
rect 3 -22 7 -18
rect 49 -5 53 -1
rect 7 -49 11 -45
rect 39 -29 43 -25
rect 61 -29 65 -25
rect 38 -37 42 -33
rect 46 -37 50 -33
rect 62 -37 66 -33
rect 78 -22 82 -18
rect 54 -49 58 -45
rect 39 -69 43 -65
rect 69 -69 73 -65
<< metal2 >>
rect 39 15 65 19
rect 49 -1 53 15
rect 13 -5 14 -1
rect 18 -5 49 -1
rect 7 -22 78 -18
rect 43 -29 61 -25
rect 42 -37 46 -33
rect 50 -37 62 -33
rect 11 -49 54 -45
rect 39 -65 43 -49
rect 43 -69 69 -65
<< labels >>
rlabel metal1 13 -3 13 -3 1 vdd
rlabel metal1 71 -27 71 -27 1 br
rlabel metal1 33 -27 33 -27 1 bl
rlabel polysilicon 13 -28 13 -28 1 din
rlabel metal1 17 -29 17 -29 1 din_bar
rlabel metal1 48 -24 48 -24 1 we_bar
rlabel polysilicon 52 -24 52 -24 1 we
rlabel metal1 37 -67 37 -67 1 gnd
<< end >>
