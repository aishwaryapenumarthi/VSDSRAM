magic
tech scmos
timestamp 1599152182
<< nwell >>
rect -8 37 35 58
rect -95 -14 -14 32
rect 41 -7 93 41
rect -5 -74 29 -29
<< ntransistor >>
rect 4 16 6 24
rect 22 16 24 24
rect 7 2 11 4
rect 17 2 21 4
rect -84 -33 -82 -29
rect -65 -34 -61 -32
rect 80 -17 82 -13
rect 50 -20 54 -18
rect 61 -20 65 -18
rect -45 -36 -43 -32
rect -27 -34 -23 -32
rect -65 -50 -61 -48
rect -27 -50 -23 -48
<< ptransistor >>
rect 4 43 6 47
rect 22 43 24 47
rect -67 14 -59 16
rect -29 14 -21 16
rect 55 19 57 30
rect 50 4 54 6
rect 58 4 66 6
rect -84 -7 -82 1
rect -67 -2 -59 0
rect -45 -7 -43 1
rect -29 -2 -21 0
rect 80 -1 82 7
rect 11 -41 13 -37
rect 3 -55 7 -53
rect 17 -55 21 -53
<< ndiffusion >>
rect -2 22 4 24
rect -2 18 -1 22
rect 3 18 4 22
rect -2 16 4 18
rect 6 22 12 24
rect 6 18 7 22
rect 11 18 12 22
rect 6 16 12 18
rect 16 22 22 24
rect 16 18 17 22
rect 21 18 22 22
rect 16 16 22 18
rect 24 23 29 24
rect 24 19 25 23
rect 24 16 29 19
rect 7 4 11 5
rect 17 4 21 5
rect 7 1 11 2
rect 17 1 21 2
rect -85 -33 -84 -29
rect -82 -33 -81 -29
rect -65 -32 -61 -31
rect -65 -35 -61 -34
rect 50 -18 54 -17
rect 79 -17 80 -13
rect 82 -17 83 -13
rect 61 -18 65 -17
rect 50 -21 54 -20
rect 61 -21 65 -20
rect -46 -36 -45 -32
rect -43 -36 -42 -32
rect -27 -32 -23 -31
rect -27 -35 -23 -34
rect -65 -48 -61 -47
rect -27 -48 -23 -47
rect -65 -51 -61 -50
rect -27 -51 -23 -50
<< pdiffusion >>
rect -2 43 -1 47
rect 3 43 4 47
rect 6 43 7 47
rect 11 43 12 47
rect 16 43 17 47
rect 21 43 22 47
rect 24 43 25 47
rect -67 17 -65 21
rect -61 17 -59 21
rect -67 16 -59 17
rect -29 17 -27 21
rect -23 17 -21 21
rect -29 16 -21 17
rect -67 13 -59 14
rect -67 9 -65 13
rect -61 9 -59 13
rect -29 13 -21 14
rect 50 23 55 30
rect 54 19 55 23
rect 57 26 58 30
rect 57 19 62 26
rect -29 9 -27 13
rect -23 9 -21 13
rect -67 1 -65 5
rect -61 1 -59 5
rect -29 1 -27 5
rect -23 1 -21 5
rect 50 6 54 7
rect 62 7 66 11
rect 58 6 66 7
rect 50 3 54 4
rect -85 -3 -84 1
rect -89 -7 -84 -3
rect -82 -3 -77 1
rect -67 0 -59 1
rect -82 -7 -81 -3
rect -67 -3 -59 -2
rect -50 -3 -45 1
rect -67 -7 -65 -3
rect -61 -7 -59 -3
rect -46 -7 -45 -3
rect -43 -3 -42 1
rect -29 0 -21 1
rect -29 -3 -21 -2
rect -43 -7 -38 -3
rect -29 -7 -27 -3
rect -23 -7 -21 -3
rect 58 3 66 4
rect 58 -1 61 3
rect 65 -1 66 3
rect 79 3 80 7
rect 75 -1 80 3
rect 82 3 87 7
rect 82 -1 83 3
rect 7 -41 11 -37
rect 13 -41 17 -37
rect 3 -53 7 -49
rect 17 -53 21 -49
rect 3 -59 7 -55
rect 17 -59 21 -55
<< ndcontact >>
rect -1 18 3 22
rect 7 18 11 22
rect 17 18 21 22
rect 25 19 29 23
rect 7 5 11 9
rect 17 5 21 9
rect 7 -3 11 1
rect 17 -3 21 1
rect -89 -33 -85 -29
rect -81 -33 -77 -29
rect -65 -31 -61 -27
rect 50 -17 54 -13
rect 61 -17 65 -13
rect 75 -17 79 -13
rect 83 -17 87 -13
rect 50 -25 54 -21
rect 61 -25 65 -21
rect -27 -31 -23 -27
rect -65 -39 -61 -35
rect -50 -36 -46 -32
rect -42 -36 -38 -32
rect -27 -39 -23 -35
rect -65 -47 -61 -43
rect -27 -47 -23 -43
rect -65 -55 -61 -51
rect -27 -55 -23 -51
<< pdcontact >>
rect -1 43 3 47
rect 7 43 11 47
rect 17 43 21 47
rect 25 43 29 47
rect -65 17 -61 21
rect -27 17 -23 21
rect -65 9 -61 13
rect 50 19 54 23
rect 58 26 62 30
rect -27 9 -23 13
rect -65 1 -61 5
rect -27 1 -23 5
rect 50 7 54 11
rect 58 7 62 11
rect -89 -3 -85 1
rect -81 -7 -77 -3
rect -65 -7 -61 -3
rect -50 -7 -46 -3
rect -42 -3 -38 1
rect -27 -7 -23 -3
rect 50 -1 54 3
rect 61 -1 65 3
rect 75 3 79 7
rect 83 -1 87 3
rect 3 -41 7 -37
rect 17 -41 21 -37
rect 3 -49 7 -45
rect 17 -49 21 -45
rect 3 -63 7 -59
rect 17 -63 21 -59
<< psubstratepcontact >>
rect -1 28 3 32
rect 25 28 29 32
rect 50 -35 54 -31
rect 75 -35 79 -31
rect -35 -55 -31 -51
rect -65 -63 -61 -59
<< nsubstratencontact >>
rect -1 51 3 55
rect 25 51 29 55
rect -65 25 -61 29
rect -27 25 -23 29
rect 50 34 54 38
rect 58 34 62 38
rect 75 12 79 16
rect 83 12 87 16
rect -89 5 -85 9
rect -42 5 -38 9
rect 3 -71 7 -67
rect 17 -71 21 -67
<< polysilicon >>
rect 4 47 6 49
rect 22 47 24 49
rect 4 40 6 43
rect 4 38 15 40
rect 4 24 6 38
rect 22 33 24 43
rect 13 31 24 33
rect 22 24 24 31
rect 55 30 57 32
rect -70 14 -67 16
rect -59 14 -57 16
rect -31 14 -29 16
rect -21 14 -18 16
rect 55 17 57 19
rect 4 14 6 16
rect 22 14 24 16
rect -84 1 -82 3
rect -45 1 -43 3
rect 5 2 7 4
rect 11 2 17 4
rect 21 2 23 4
rect 80 7 82 9
rect 45 4 50 6
rect 54 4 58 6
rect 66 4 68 6
rect -69 -2 -67 0
rect -59 -2 -57 0
rect -31 -2 -29 0
rect -21 -2 -19 0
rect -84 -29 -82 -7
rect -45 -16 -43 -7
rect 13 -10 15 2
rect 80 -9 82 -1
rect 71 -11 82 -9
rect 80 -13 82 -11
rect -45 -18 -40 -16
rect -84 -35 -82 -33
rect -67 -34 -65 -32
rect -61 -34 -58 -32
rect -45 -32 -43 -18
rect 47 -20 50 -18
rect 54 -20 56 -18
rect 59 -20 61 -18
rect 65 -20 68 -18
rect 80 -19 82 -17
rect -30 -34 -27 -32
rect -23 -34 -21 -32
rect -45 -38 -43 -36
rect 11 -37 13 -35
rect -70 -50 -65 -48
rect -61 -50 -59 -48
rect -29 -50 -27 -48
rect -23 -50 -18 -48
rect 11 -53 13 -41
rect 1 -55 3 -53
rect 7 -55 10 -53
rect 14 -55 17 -53
rect 21 -55 23 -53
<< polycontact >>
rect 15 37 19 41
rect 9 30 13 34
rect -74 13 -70 17
rect -18 13 -14 17
rect 41 3 45 7
rect -57 -3 -53 1
rect -35 -3 -31 1
rect -88 -12 -84 -8
rect 12 -14 16 -10
rect 67 -12 71 -8
rect -58 -35 -54 -31
rect -40 -19 -36 -15
rect 43 -21 47 -17
rect 68 -21 72 -17
rect -34 -35 -30 -31
rect -74 -51 -70 -47
rect -18 -51 -14 -47
rect 10 -57 14 -53
<< metal1 >>
rect 3 51 25 55
rect -1 47 3 51
rect 25 47 29 51
rect 7 34 11 43
rect 17 41 21 43
rect 19 37 21 41
rect -65 21 -61 25
rect -27 21 -23 25
rect -1 22 3 28
rect 7 30 9 34
rect 7 29 11 30
rect 7 22 11 25
rect 17 29 21 37
rect 54 34 58 38
rect 17 22 21 25
rect 25 23 29 28
rect 58 30 62 34
rect -85 5 -82 9
rect -89 1 -85 5
rect -89 -12 -88 -8
rect -81 -17 -77 -7
rect -74 -17 -70 13
rect -65 5 -61 9
rect -43 5 -42 9
rect -42 1 -38 5
rect -27 5 -23 9
rect -81 -21 -70 -17
rect -81 -29 -77 -21
rect -89 -39 -85 -33
rect -74 -47 -70 -21
rect -65 -15 -61 -7
rect -57 -15 -53 -3
rect -65 -19 -60 -15
rect -65 -27 -61 -19
rect -50 -27 -46 -7
rect -35 -15 -31 -3
rect -36 -19 -35 -15
rect -27 -23 -23 -7
rect -50 -32 -46 -31
rect -18 -8 -14 13
rect -1 10 3 18
rect 7 9 11 10
rect 17 9 21 10
rect 25 10 29 19
rect 50 16 54 19
rect 50 12 62 16
rect 50 11 54 12
rect 58 11 62 12
rect 79 12 83 16
rect 75 7 79 12
rect 41 -1 50 3
rect -65 -43 -61 -39
rect -42 -39 -38 -36
rect -27 -43 -23 -39
rect -18 -47 -14 -12
rect -1 -14 12 -10
rect 16 -14 29 -10
rect 50 -13 54 -1
rect 61 -8 65 -1
rect 83 -8 87 -1
rect 61 -12 67 -8
rect 83 -12 88 -8
rect 61 -13 65 -12
rect 83 -13 87 -12
rect 50 -31 54 -25
rect 61 -31 65 -25
rect 68 -24 72 -21
rect 75 -31 79 -17
rect 3 -37 7 -31
rect 3 -45 7 -41
rect 54 -35 75 -31
rect 17 -45 21 -41
rect -31 -55 -27 -51
rect -65 -59 -61 -55
rect -27 -59 -23 -55
rect -61 -63 -57 -59
rect 10 -61 14 -57
rect 3 -67 7 -63
rect 17 -67 21 -63
rect 7 -71 17 -67
<< m2contact >>
rect -61 25 -57 29
rect -31 25 -27 29
rect 7 25 11 29
rect 17 25 21 29
rect -82 5 -78 9
rect -93 -12 -89 -8
rect -47 5 -43 9
rect -89 -43 -85 -39
rect -57 -19 -53 -15
rect -35 -19 -31 -15
rect -27 -27 -23 -23
rect -58 -31 -54 -27
rect -50 -31 -46 -27
rect -34 -31 -30 -27
rect -1 6 3 10
rect 7 10 11 14
rect 17 10 21 14
rect 25 6 29 10
rect 7 -7 11 -3
rect 17 -7 21 -3
rect -18 -12 -14 -8
rect -42 -43 -38 -39
rect 39 -21 43 -17
rect 68 -28 72 -24
rect 17 -37 21 -33
rect -57 -63 -53 -59
rect -27 -63 -23 -59
<< metal2 >>
rect -57 25 -31 29
rect -47 9 -43 25
rect 7 14 11 25
rect 17 14 21 25
rect 25 10 29 14
rect -83 5 -82 9
rect -78 5 -47 9
rect -89 -12 -18 -8
rect -1 -14 3 6
rect 7 -15 11 -7
rect -53 -19 -35 -15
rect 17 -17 21 -7
rect 25 -14 29 6
rect 17 -21 39 -17
rect 17 -23 21 -21
rect -23 -27 21 -23
rect -54 -31 -50 -27
rect -46 -31 -34 -27
rect 17 -33 21 -27
rect 43 -28 68 -24
rect -85 -43 -42 -39
rect -57 -59 -53 -43
rect -53 -63 -27 -59
<< m3contact >>
rect -65 -19 -60 -15
rect 7 -20 11 -15
rect 3 -36 7 -31
rect 38 -28 43 -24
<< metal3 >>
rect -60 -19 7 -15
rect 3 -24 7 -19
rect 3 -28 38 -24
rect 3 -31 7 -28
<< labels >>
rlabel metal1 -83 7 -83 7 1 vdd
rlabel polysilicon -83 -18 -83 -18 1 din
rlabel metal1 -79 -19 -79 -19 1 din_bar
rlabel metal1 -59 -61 -59 -61 1 gnd
rlabel metal1 -25 -17 -25 -17 1 br
rlabel polysilicon -44 -14 -44 -14 1 we
rlabel metal1 -48 -14 -48 -14 1 we_bar
rlabel metal1 -63 -17 -63 -17 1 bl
rlabel metal1 9 36 9 36 1 q
rlabel metal1 1 14 1 14 1 gnd
rlabel m2contact 9 -4 9 -4 1 bl
rlabel m2contact 19 -4 19 -4 1 br
rlabel metal1 27 14 27 14 1 gnd
rlabel metal1 19 35 19 35 1 qb
rlabel metal1 15 53 15 53 5 vdd
rlabel metal1 18 -12 18 -12 1 wl
rlabel m2contact 19 -35 19 -35 1 br
rlabel metal1 12 -59 12 -59 5 pre
rlabel metal1 12 -69 12 -69 5 vdd
rlabel metal1 5 -35 5 -35 5 bl
rlabel metal1 57 -33 57 -33 1 gnd
rlabel metal1 88 -12 88 -8 7 dout
rlabel metal1 81 14 81 14 1 vdd
rlabel metal1 64 -10 64 -10 1 amp_out
rlabel metal1 56 36 56 36 5 vdd
rlabel polysilicon 55 32 57 32 1 sen
<< end >>
