* SPICE3 file created from Integrated.ext - technology: scmos
.include osu018.lib
.option scale=0.1u

M1000 q wl bl gnd nfet w=4 l=2
+  ad=68 pd=46 as=40 ps=36
M1001 dout amp_out vdd vdd pfet w=8 l=2
+  ad=40 pd=26 as=363 ps=248
M1002 a_41_3# br gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=228 ps=180
M1003 amp_out bl gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 br pre bl vdd pfet w=4 l=2
+  ad=104 pd=74 as=104 ps=74
M1005 q qb vdd vdd pfet w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1006 vdd din_bar a_n67_0# vdd pfet w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1007 gnd we we_bar gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1008 br we_bar a_n27_n48# gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1009 vdd we we_bar vdd pfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1010 din_bar din vdd vdd pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1011 a_n29_0# we br vdd pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1012 a_n65_n48# din_bar gnd gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1013 vdd sen a_50_6# vdd pfet w=11 l=2
+  ad=0 pd=0 as=115 ps=76
M1014 a_50_6# a_41_3# a_41_3# vdd pfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1015 dout amp_out gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1016 br pre vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 gnd q qb gnd nfet w=8 l=2
+  ad=0 pd=0 as=68 ps=46
M1018 qb wl br gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 vdd din a_n29_0# vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 a_50_6# a_41_3# amp_out vdd pfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1021 vdd q qb vdd pfet w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1022 bl we_bar a_n65_n48# gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 a_n27_n48# din gnd gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 bl pre vdd vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 din_bar din gnd gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1026 a_n67_0# we bl vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 q qb gnd gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 br a_n29_0# 0.04fF
C1 bl amp_out 0.05fF
C2 a_n27_n48# br 0.04fF
C3 a_n67_0# din_bar 0.10fF
C4 a_n65_n48# din_bar 0.10fF
C5 vdd we 0.41fF
C6 amp_out a_50_6# 0.01fF
C7 vdd bl 0.09fF
C8 din din_bar 0.11fF
C9 br din 0.28fF
C10 vdd a_50_6# 0.08fF
C11 a_41_3# a_50_6# 0.04fF
C12 vdd pre 0.35fF
C13 bl wl 0.08fF
C14 we_bar din 0.03fF
C15 vdd a_n29_0# 0.06fF
C16 bl we 0.31fF
C17 vdd a_n67_0# 0.09fF
C18 br we_bar 0.05fF
C19 vdd din 0.40fF
C20 qb br 0.04fF
C21 vdd dout 0.03fF
C22 vdd din_bar 0.31fF
C23 bl a_n67_0# 0.04fF
C24 q qb 0.59fF
C25 vdd br 0.09fF
C26 bl a_n65_n48# 0.04fF
C27 vdd sen 0.05fF
C28 we din 0.47fF
C29 bl din 0.11fF
C30 q vdd 0.17fF
C31 vdd we_bar 0.03fF
C32 br wl 0.08fF
C33 bl din_bar 0.23fF
C34 qb vdd 0.27fF
C35 vdd amp_out 0.09fF
C36 amp_out a_41_3# 0.12fF
C37 br we 0.16fF
C38 bl br 0.49fF
C39 a_n29_0# din 0.10fF
C40 a_n27_n48# din 0.10fF
C41 vdd a_41_3# 0.20fF
C42 we_bar we 0.28fF
C43 q bl 0.04fF
C44 bl we_bar 0.06fF
C45 bl gnd 0.32fF
C46 a_n27_n48# gnd 0.03fF
C47 a_n65_n48# gnd 0.03fF
C48 dout gnd 0.04fF
C49 br gnd 0.10fF
C50 we_bar gnd 0.36fF
C51 amp_out gnd 0.22fF
C52 a_41_3# gnd 0.05fF
C53 wl gnd 0.31fF
C54 we gnd 0.29fF
C55 a_n29_0# gnd 0.00fF
C56 a_n67_0# gnd 0.00fF
C57 din gnd 0.42fF
C58 din_bar gnd 0.33fF
C59 q gnd 0.52fF
C60 qb gnd 0.46fF
C61 vdd gnd 5.44fF


*voltages


v1 vdd gnd  dc 1.8V

v2 wl gnd pulse(0V 1.8V 0ns 1ns 1ns 50ns 100ns)

v3 pre gnd pulse(1.8V 0V 50ns 1ns 1ns 50ns 100ns)

v6 we gnd pulse(1.8V 0V 0ns 1ns 1ns 50ns 100ns)

v7 sen gnd pulse(0V 1.8V 50ns 1ns 1ns 50ns 100ns)

v8 din gnd pulse(0V 1.8V 0ns 1ns 1ns 10ns 20ns)

.tran 10e-12 200e-09 1e-09

.control
run

plot v(wl)+12 v(we)+10 v(din)+8 v(sen)+6 v(pre)+4  v(dout)

plot v(bl)+2 v(br)


.endc
.end
