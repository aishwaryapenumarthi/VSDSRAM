* SPICE3 file created from precharge.ext - technology: scmos

.option scale=0.1u
.include osu018.lib

M1000 vdd pre br vdd pfet w=4 l=2
+  ad=64 pd=48 as=64 ps=48
M1001 bl pre br vdd pfet w=4 l=2
+  ad=64 pd=48 as=0 ps=0
M1002 vdd pre bl vdd pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0

v1  vdd gnd 1.8V
v2  pre gnd pulse(0 1.8V 50ps 10ps 10ps 40ns 80ns)
.tran 10e-09 100e-09 0e-09

* Control Statements 
.control
run

plot v(pre)+6 v(bl)+3 v(br)

.endc
.end
