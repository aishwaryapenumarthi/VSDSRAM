magic
tech sample_6m
timestamp 1598000048
<< nwell >>
rect -58 -35 -20 34
rect -6 -36 23 -1
<< ntransistor >>
rect -50 -53 -46 -51
rect -32 -53 -28 -51
rect 7 -50 9 -46
<< ptransistor >>
rect -41 -2 -39 12
rect -49 -21 -45 -19
rect -35 -21 -25 -19
rect 7 -31 9 -21
<< ndiffusion >>
rect -50 -51 -46 -49
rect -32 -51 -28 -49
rect -50 -55 -46 -53
rect -32 -55 -28 -53
rect 4 -50 7 -46
rect 9 -50 12 -46
<< pdiffusion >>
rect -51 5 -41 12
rect -51 0 -50 5
rect -45 0 -41 5
rect -51 -2 -41 0
rect -39 10 -29 12
rect -39 5 -35 10
rect -30 5 -29 10
rect -39 -2 -29 5
rect -49 -19 -45 -16
rect -35 -16 -34 -11
rect -29 -16 -25 -11
rect -35 -19 -25 -16
rect -49 -24 -45 -21
rect -35 -24 -25 -21
rect -35 -29 -32 -24
rect -27 -29 -25 -24
rect 4 -26 7 -21
rect -1 -31 7 -26
rect 9 -26 17 -21
rect 9 -31 12 -26
<< ndcontact >>
rect -50 -49 -45 -44
rect -32 -49 -27 -44
rect -1 -51 4 -46
rect 12 -50 17 -45
rect -50 -60 -45 -55
rect -32 -60 -27 -55
<< pdcontact >>
rect -50 0 -45 5
rect -35 5 -30 10
rect -50 -16 -45 -11
rect -34 -16 -29 -11
rect -50 -29 -45 -24
rect -32 -29 -27 -24
rect -1 -26 4 -21
rect 12 -31 17 -26
<< psubstratepcontact >>
rect -1 -66 4 -61
rect 14 -66 19 -61
rect -50 -75 -45 -70
rect -32 -75 -27 -70
<< nsubstratencontact >>
rect -51 24 -46 29
rect -35 24 -30 29
rect -1 -11 4 -6
rect 14 -11 19 -6
<< polysilicon >>
rect -41 12 -39 16
rect -41 -5 -39 -2
rect -52 -21 -49 -19
rect -45 -21 -35 -19
rect -25 -21 -22 -19
rect 7 -21 9 -18
rect 7 -38 9 -31
rect 8 -43 9 -38
rect 7 -46 9 -43
rect -54 -53 -50 -51
rect -46 -53 -43 -51
rect -35 -53 -32 -51
rect -28 -53 -24 -51
rect 7 -53 9 -50
<< polycontact >>
rect -43 16 -38 21
rect -57 -24 -52 -19
rect 3 -43 8 -38
rect -59 -54 -54 -49
rect -24 -54 -19 -49
<< metal1 >>
rect -46 24 -35 29
rect -44 16 -43 21
rect -35 10 -30 24
rect -50 -11 -45 0
rect 4 -11 14 -6
rect -45 -16 -34 -11
rect -1 -21 4 -11
rect -57 -29 -50 -24
rect -50 -44 -45 -29
rect -32 -38 -27 -29
rect 12 -38 17 -31
rect -32 -43 3 -38
rect 12 -42 19 -38
rect -32 -44 -27 -43
rect 12 -45 17 -42
rect -62 -54 -59 -49
rect -19 -54 -16 -49
rect -50 -70 -45 -60
rect -32 -70 -27 -60
rect -1 -61 4 -51
rect 4 -66 14 -61
rect -45 -75 -32 -70
<< labels >>
rlabel metal1 -44 16 -44 21 1 sen
rlabel metal1 -16 -54 -16 -49 1 bl
rlabel metal1 -62 -54 -62 -49 3 br
rlabel metal1 9 -64 9 -64 1 gnd
rlabel metal1 -39 -73 -39 -73 1 gnd
rlabel metal1 -40 27 -40 27 1 vdd
rlabel metal1 9 -8 9 -8 1 vdd
rlabel metal1 19 -42 19 -38 7 dout
<< end >>
