* SPICE3 file created from writedriver.ext - technology: sample_6m

.include osu018.lib
.option scale=0.09u

M1000 gnd we a_4_n29# gnd nmos w=5 l=2
+  ad=150 pd=100 as=40 ps=26
M1001 a_5_0# we bl vdd pmos w=10 l=2
+  ad=140 pd=68 as=70 ps=34
M1002 vdd we a_4_n29# vdd pmos w=10 l=2
+  ad=300 pd=140 as=80 ps=36
M1003 vdd din a_88_2# vdd pmos w=10 l=2
+  ad=0 pd=0 as=140 ps=68
M1004 a_88_2# we br vdd pmos w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1005 br a_4_n29# a_91_n46# gnd nmos w=5 l=2
+  ad=35 pd=24 as=70 ps=48
M1006 a_n37_n21# din gnd gnd nmos w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1007 a_91_n46# din gnd gnd nmos w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 bl a_4_n29# a_7_n48# gnd nmos w=5 l=2
+  ad=35 pd=24 as=70 ps=48
M1009 a_7_n48# a_n37_n21# gnd gnd nmos w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 vdd a_n37_n21# a_5_0# vdd pmos w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_n37_n21# din vdd vdd pmos w=10 l=2
+  ad=80 pd=36 as=0 ps=0



v1  din gnd pulse(0 1.8V 0 100ps 100ps 10ns 20ns)
v2  vdd gnd 1.8v
v3  we gnd pulse(0 1.8V 0 100ps 100ps 50ns 100ns)
.tran 10e-09 100e-09 0e-09
.control
run

plot v(we)+9 v(din)+6 v(bl)+3 v(br)

.endc
.end
