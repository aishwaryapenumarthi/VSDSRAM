* SPICE3 file created from new_dflipflop.ext - technology: scmos

.option scale=0.1u
.include osu018.lib


M1000 S d_bar net2 gnd nfet w=4 l=2
+  ad=40 pd=36 as=20 ps=18
M1001 gnd d d_bar gnd nfet w=4 l=2
+  ad=100 pd=90 as=20 ps=18
M1002 gnd clk P gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1003 gnd qb U gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1004 gnd q T gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1005 net1 d vdd vdd pfet w=7 l=2
+  ad=75 pd=50 as=355 ps=232
M1006 net2 d_bar vdd vdd pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1007 vdd d d_bar vdd pfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1008 gnd clk S gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 P d net1 gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1010 U net1 q gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1011 T net2 qb gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1012 qb net2 vdd vdd pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1013 q net1 vdd vdd pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1014 net2 clk vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 net1 clk vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 q qb vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 qb q vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 clk net1 0.08fF
C1 net1 d 0.08fF
C2 qb net1 0.02fF
C3 clk d_bar 0.02fF
C4 S net2 0.04fF
C5 d_bar d 0.05fF
C6 clk vdd 0.21fF
C7 net1 P 0.04fF
C8 net2 d_bar 0.05fF
C9 d vdd 0.22fF
C10 qb vdd 0.23fF
C11 q qb 0.18fF
C12 net2 vdd 0.24fF
C13 U vdd 0.03fF
C14 q net2 0.02fF
C15 P vdd 0.03fF
C16 net1 vdd 0.31fF
C17 q U 0.04fF
C18 q net1 0.03fF
C19 d_bar vdd 0.19fF
C20 T qb 0.04fF
C21 q vdd 0.31fF
C22 clk d 0.01fF
C23 clk net2 0.08fF
C24 qb net2 0.03fF
C25 T gnd 0.03fF
C26 U gnd 0.03fF
C27 qb gnd 0.76fF
C28 q gnd 0.95fF
C29 S gnd 0.03fF
C30 P gnd 0.03fF
C31 clk gnd 0.25fF
C32 net2 gnd 0.40fF
C33 net1 gnd 0.38fF
C34 d_bar gnd 0.39fF
C35 d gnd 0.60fF
C36 vdd gnd 3.91fF


v3 vdd gnd  dc 1.8V
v2  d gnd pulse(0 1.8V 0 10ps 10ps 10ns 20ns)
v1  clk gnd pulse(0 1.8V 0 10ps 10ps 50ns 100ns)

.tran 10e-09 100e-09 0e-09

* Control Statements 
.control
run
plot v(clk)+6 v(d)+4 v(q)+2 v(qb)
.endc
.end
