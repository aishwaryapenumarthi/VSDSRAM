magic
tech sample_6m
timestamp 1598115420
<< nwell >>
rect -4 -5 22 23
rect 37 -5 63 23
<< ntransistor >>
rect -35 -10 -33 -6
rect 8 -20 10 -12
rect 91 -11 93 -7
rect 49 -21 51 -13
<< ptransistor >>
rect 8 1 10 5
rect 49 1 51 5
<< ndiffusion >>
rect -37 -10 -35 -6
rect -33 -10 -31 -6
rect 1 -13 8 -12
rect 6 -18 8 -13
rect 1 -20 8 -18
rect 10 -14 17 -12
rect 89 -11 91 -7
rect 93 -11 95 -7
rect 10 -19 12 -14
rect 10 -20 17 -19
rect 42 -15 49 -13
rect 47 -20 49 -15
rect 42 -21 49 -20
rect 51 -14 58 -13
rect 51 -19 53 -14
rect 51 -21 58 -19
<< pdiffusion >>
rect 6 1 8 5
rect 10 1 12 5
rect 47 1 49 5
rect 51 1 53 5
<< ndcontact >>
rect -42 -11 -37 -6
rect -31 -11 -26 -6
rect 1 -18 6 -13
rect 84 -12 89 -7
rect 12 -19 17 -14
rect 42 -20 47 -15
rect 95 -12 100 -7
rect 53 -19 58 -14
<< pdcontact >>
rect 1 0 6 5
rect 12 1 17 6
rect 42 1 47 6
rect 53 0 58 5
<< psubstratepcontact >>
rect 1 -35 6 -30
rect 12 -35 17 -30
rect 42 -36 47 -31
rect 53 -36 58 -31
<< nsubstratencontact >>
rect 1 16 6 21
rect 12 16 17 21
rect 42 16 47 21
rect 53 16 58 21
<< polysilicon >>
rect -35 36 93 38
rect -35 -6 -33 36
rect 8 28 67 30
rect 8 5 10 28
rect 49 5 51 8
rect -35 -13 -33 -10
rect -8 -40 -6 -11
rect 8 -12 10 1
rect 49 -13 51 1
rect 65 -7 67 28
rect 91 -7 93 36
rect 8 -23 10 -20
rect 91 -14 93 -11
rect 49 -25 51 -21
rect 49 -27 68 -25
rect 66 -40 68 -27
rect -8 -42 68 -40
<< polycontact >>
rect -10 -11 -5 -6
rect 64 -12 69 -7
<< metal1 >>
rect 6 16 12 21
rect 12 6 17 16
rect 47 16 53 21
rect 42 6 47 16
rect 1 -6 6 0
rect -45 -11 -42 -6
rect -26 -11 -10 -6
rect -5 -11 6 -6
rect 1 -13 6 -11
rect 53 -7 58 0
rect 53 -12 64 -7
rect 69 -12 84 -7
rect 100 -12 104 -7
rect 53 -14 58 -12
rect 12 -30 17 -19
rect 6 -35 12 -30
rect 42 -31 47 -20
rect 47 -36 53 -31
<< labels >>
rlabel metal1 -45 -11 -45 -6 3 bl
rlabel metal1 104 -12 104 -7 7 br
rlabel metal1 60 -9 60 -9 1 qb
rlabel metal1 4 -8 4 -8 1 q
rlabel metal1 11 19 11 19 1 vdd
rlabel metal1 50 18 50 18 1 vdd
rlabel metal1 9 -33 9 -33 1 gnd
rlabel metal1 51 -34 51 -34 1 gnd
rlabel polysilicon 32 37 32 37 5 wl
<< end >>
