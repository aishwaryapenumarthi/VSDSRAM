magic
tech scmos
timestamp 1598304036
<< nwell >>
rect -7 -2 17 20
rect 25 -2 49 20
<< ntransistor >>
rect -26 -7 -24 -3
rect 69 -7 71 -3
rect 4 -16 6 -8
rect 36 -16 38 -8
<< ptransistor >>
rect 4 4 6 8
rect 36 4 38 8
<< ndiffusion >>
rect -27 -7 -26 -3
rect -24 -7 -23 -3
rect 68 -7 69 -3
rect 71 -7 72 -3
rect 3 -12 4 -8
rect -1 -16 4 -12
rect 6 -12 11 -8
rect 6 -16 7 -12
rect 31 -12 36 -8
rect 35 -16 36 -12
rect 38 -12 39 -8
rect 38 -16 43 -12
<< pdiffusion >>
rect 3 4 4 8
rect 6 4 7 8
rect 35 4 36 8
rect 38 4 39 8
<< ndcontact >>
rect -31 -7 -27 -3
rect -23 -7 -19 -3
rect 64 -7 68 -3
rect 72 -7 76 -3
rect -1 -12 3 -8
rect 7 -16 11 -12
rect 31 -16 35 -12
rect 39 -12 43 -8
<< pdcontact >>
rect -1 4 3 8
rect 7 4 11 8
rect 31 4 35 8
rect 39 4 43 8
<< psubstratepcontact >>
rect -1 -25 3 -21
rect 7 -25 11 -21
rect 31 -25 35 -21
rect 40 -25 44 -21
<< nsubstratencontact >>
rect -2 13 2 17
rect 7 13 11 17
rect 31 13 35 17
rect 40 13 44 17
<< polysilicon >>
rect -26 26 71 28
rect -26 -3 -24 26
rect 4 21 53 23
rect 4 8 6 21
rect 36 8 38 10
rect -26 -10 -24 -7
rect -10 -33 -8 -7
rect 4 -8 6 4
rect 36 -8 38 4
rect 51 -3 53 21
rect 69 -3 71 26
rect 69 -10 71 -7
rect 4 -18 6 -16
rect 36 -33 38 -16
rect -10 -35 38 -33
<< polycontact >>
rect -11 -7 -7 -3
rect 50 -7 54 -3
<< metal1 >>
rect 2 13 7 17
rect 7 8 11 13
rect 35 13 40 17
rect 31 8 35 13
rect -1 -3 3 4
rect -32 -7 -31 -3
rect -19 -7 -11 -3
rect -7 -7 3 -3
rect -1 -8 3 -7
rect 39 -3 43 4
rect 39 -7 50 -3
rect 54 -7 64 -3
rect 76 -7 77 -3
rect 39 -8 43 -7
rect 7 -21 11 -16
rect 3 -25 7 -21
rect 31 -21 35 -16
rect 35 -25 40 -21
<< labels >>
rlabel metal1 1 -5 1 -5 1 q
rlabel metal1 41 -5 41 -5 1 qb
rlabel metal1 77 -7 77 -3 7 br
rlabel metal1 -32 -7 -32 -3 3 bl
rlabel metal1 5 -23 5 -23 1 gnd
rlabel polysilicon 30 27 30 27 5 wl
rlabel metal1 3 15 3 15 1 vdd
rlabel metal1 37 15 37 15 1 vdd
rlabel metal1 39 -23 39 -23 1 gnd
<< end >>
