magic
tech sample_6m
timestamp 1598192121
<< nwell >>
rect -50 -24 -21 9
rect 0 -14 23 44
rect 33 3 62 36
<< ntransistor >>
rect 46 -9 48 -5
rect 7 -29 12 -27
rect -36 -36 -34 -32
rect 7 -50 12 -48
<< ptransistor >>
rect 5 18 14 20
rect 46 9 48 19
rect 5 -2 14 0
rect -36 -18 -34 -8
<< ndiffusion >>
rect 43 -9 46 -5
rect 48 -9 51 -5
rect 7 -21 12 -20
rect 7 -27 12 -26
rect 7 -30 12 -29
rect -39 -36 -36 -32
rect -34 -36 -31 -32
rect 7 -36 12 -35
rect 7 -42 12 -41
rect 7 -48 12 -47
rect 7 -52 12 -50
<< pdiffusion >>
rect 5 26 14 27
rect 5 21 7 26
rect 12 21 14 26
rect 5 20 14 21
rect 5 17 14 18
rect 5 12 7 17
rect 12 12 14 17
rect 5 11 14 12
rect 38 14 46 19
rect 43 9 46 14
rect 48 14 51 19
rect 48 9 56 14
rect 5 6 14 7
rect 5 1 7 6
rect 12 1 14 6
rect 5 0 14 1
rect 5 -3 14 -2
rect 5 -8 7 -3
rect 12 -8 14 -3
rect -39 -13 -36 -8
rect -44 -18 -36 -13
rect -34 -13 -26 -8
rect 5 -9 14 -8
rect -34 -18 -31 -13
<< ndcontact >>
rect 38 -9 43 -4
rect 51 -10 56 -5
rect 7 -26 12 -21
rect -44 -37 -39 -32
rect -31 -36 -26 -31
rect 7 -35 12 -30
rect 7 -47 12 -42
rect 7 -57 12 -52
<< pdcontact >>
rect 7 21 12 26
rect 7 12 12 17
rect 38 9 43 14
rect 51 14 56 19
rect 7 1 12 6
rect 7 -8 12 -3
rect -44 -13 -39 -8
rect -31 -18 -26 -13
<< psubstratepcontact >>
rect 38 -25 43 -20
rect 51 -25 56 -20
rect -44 -52 -39 -47
rect -31 -52 -26 -47
rect 7 -72 12 -67
rect 17 -72 22 -67
<< nsubstratencontact >>
rect 7 37 12 42
rect 16 37 21 42
rect 39 29 44 34
rect 51 29 56 34
rect -44 2 -39 7
rect -32 2 -27 7
<< polysilicon >>
rect -2 18 5 20
rect 14 18 17 20
rect 46 19 48 22
rect 2 -2 5 0
rect 14 -2 25 0
rect 46 0 48 9
rect 46 -2 59 0
rect -36 -8 -34 -5
rect 46 -5 48 -2
rect 46 -12 48 -9
rect -36 -32 -34 -18
rect 57 -27 59 -2
rect 4 -29 7 -27
rect 12 -29 59 -27
rect -36 -39 -34 -36
rect 3 -50 7 -48
rect 12 -50 15 -48
<< polycontact >>
rect -7 16 -2 21
rect 25 -3 30 2
rect -2 -51 3 -46
<< metal1 >>
rect 12 37 16 42
rect 21 37 22 42
rect 7 26 12 37
rect 44 29 51 34
rect -19 16 -7 21
rect 51 19 56 29
rect -39 2 -32 7
rect -44 -8 -39 2
rect -31 -25 -26 -18
rect -19 -25 -14 16
rect 7 6 12 12
rect 38 2 43 9
rect 30 -3 43 2
rect -31 -30 -14 -25
rect 7 -15 12 -8
rect 38 -4 43 -3
rect 7 -19 13 -15
rect 7 -21 12 -19
rect 51 -20 56 -10
rect 43 -25 51 -20
rect -31 -31 -26 -30
rect -44 -47 -39 -37
rect -19 -46 -14 -30
rect 7 -42 12 -35
rect -39 -52 -31 -47
rect -19 -51 -2 -46
rect 7 -52 12 -51
rect 7 -67 12 -57
rect 12 -72 17 -67
<< labels >>
rlabel metal1 13 -19 13 -15 1 out
rlabel metal1 14 -69 14 -69 1 gnd
rlabel metal1 13 40 13 40 5 vdd
rlabel polysilicon -35 -27 -35 -27 3 in
rlabel metal1 -35 5 -35 5 5 vdd
rlabel metal1 -35 -50 -35 -50 3 gnd
rlabel metal1 47 32 47 32 5 vdd
rlabel metal1 47 -22 47 -22 7 gnd
rlabel polysilicon 57 -1 57 -1 7 en
<< end >>
