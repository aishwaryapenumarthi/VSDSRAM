magic
tech scmos
timestamp 1598302308
<< nwell >>
rect -2 -23 24 20
<< ptransistor >>
rect 4 0 8 2
rect 14 0 18 2
rect 10 -17 12 -13
<< pdiffusion >>
rect 4 2 8 5
rect 14 2 18 5
rect 4 -3 8 0
rect 14 -3 18 0
rect 8 -17 10 -13
rect 12 -17 14 -13
<< pdcontact >>
rect 4 5 8 9
rect 14 5 18 9
rect 4 -7 8 -3
rect 14 -7 18 -3
rect 4 -17 8 -13
rect 14 -17 18 -13
<< nsubstratencontact >>
rect 4 13 8 17
rect 14 13 18 17
<< polysilicon >>
rect 2 0 4 2
rect 8 0 14 2
rect 18 0 20 2
rect 10 -13 12 0
rect 10 -19 12 -17
<< metal1 >>
rect 8 13 14 17
rect 4 9 8 13
rect 14 9 18 13
rect 4 -13 8 -7
rect 4 -18 8 -17
rect 14 -13 18 -7
rect 14 -18 18 -17
<< labels >>
rlabel polysilicon 11 1 11 1 1 pre
rlabel metal1 11 15 11 15 1 vdd
rlabel metal1 4 -18 8 -18 1 bl
rlabel metal1 14 -18 18 -18 1 br
<< end >>
