magic
tech scmos
timestamp 1599154764
<< nwell >>
rect -26 -23 26 25
<< ntransistor >>
rect 13 -33 15 -29
rect -17 -36 -13 -34
rect -6 -36 -2 -34
<< ptransistor >>
rect -12 3 -10 14
rect -17 -12 -13 -10
rect -9 -12 -1 -10
rect 13 -17 15 -9
<< ndiffusion >>
rect -17 -34 -13 -33
rect 12 -33 13 -29
rect 15 -33 16 -29
rect -6 -34 -2 -33
rect -17 -37 -13 -36
rect -6 -37 -2 -36
<< pdiffusion >>
rect -17 7 -12 14
rect -13 3 -12 7
rect -10 10 -9 14
rect -10 3 -5 10
rect -17 -10 -13 -9
rect -5 -9 -1 -5
rect -9 -10 -1 -9
rect -17 -13 -13 -12
rect -9 -13 -1 -12
rect -9 -17 -6 -13
rect -2 -17 -1 -13
rect 12 -13 13 -9
rect 8 -17 13 -13
rect 15 -13 20 -9
rect 15 -17 16 -13
<< ndcontact >>
rect -17 -33 -13 -29
rect -6 -33 -2 -29
rect 8 -33 12 -29
rect 16 -33 20 -29
rect -17 -41 -13 -37
rect -6 -41 -2 -37
<< pdcontact >>
rect -17 3 -13 7
rect -9 10 -5 14
rect -17 -9 -13 -5
rect -9 -9 -5 -5
rect -17 -17 -13 -13
rect -6 -17 -2 -13
rect 8 -13 12 -9
rect 16 -17 20 -13
<< psubstratepcontact >>
rect -17 -51 -13 -47
rect 8 -51 12 -47
<< nsubstratencontact >>
rect -17 18 -13 22
rect -9 18 -5 22
rect 8 -4 12 0
rect 16 -4 20 0
<< polysilicon >>
rect -12 14 -10 16
rect -12 1 -10 3
rect 13 -9 15 -7
rect -22 -12 -17 -10
rect -13 -12 -9 -10
rect -1 -12 1 -10
rect 13 -25 15 -17
rect 4 -27 15 -25
rect 13 -29 15 -27
rect -20 -36 -17 -34
rect -13 -36 -11 -34
rect -8 -36 -6 -34
rect -2 -36 1 -34
rect 13 -35 15 -33
<< polycontact >>
rect -26 -13 -22 -9
rect 0 -28 4 -24
rect -24 -37 -20 -33
rect 1 -37 5 -33
<< metal1 >>
rect -13 18 -9 22
rect -9 14 -5 18
rect -17 0 -13 3
rect -17 -4 -5 0
rect -17 -5 -13 -4
rect -9 -5 -5 -4
rect 12 -4 16 0
rect 8 -9 12 -4
rect -26 -17 -17 -13
rect -17 -29 -13 -17
rect -6 -24 -2 -17
rect 16 -24 20 -17
rect -6 -28 0 -24
rect 16 -28 21 -24
rect -6 -29 -2 -28
rect 16 -29 20 -28
rect -26 -37 -24 -33
rect -17 -47 -13 -41
rect -6 -47 -2 -41
rect 1 -40 5 -37
rect 8 -47 12 -33
rect -13 -51 8 -47
<< m2contact >>
rect 1 -44 5 -40
<< metal2 >>
rect -26 -44 1 -40
<< labels >>
rlabel metal1 -10 -49 -10 -49 1 gnd
rlabel metal1 21 -28 21 -24 7 dout
rlabel metal1 14 -2 14 -2 1 vdd
rlabel metal1 -3 -26 -3 -26 1 amp_out
rlabel metal1 -11 20 -11 20 5 vdd
rlabel polysilicon -12 16 -10 16 1 sen
rlabel metal2 -23 -42 -23 -42 3 bl
rlabel metal1 -25 -35 -25 -35 3 br
<< end >>
