magic
tech scmos
timestamp 1598399373
<< nwell >>
rect -65 -9 -41 17
rect -29 -3 -9 43
rect 46 12 70 38
rect 110 -3 130 43
rect 48 -88 72 -51
rect 29 -119 53 -98
rect 59 -119 83 -98
rect 6 -188 30 -162
rect 36 -199 74 -147
<< ntransistor >>
rect 57 2 59 6
rect -54 -19 -52 -15
rect -21 -16 -17 -14
rect 118 -16 122 -14
rect -21 -32 -17 -30
rect 118 -32 122 -30
rect 16 -125 18 -121
rect 94 -124 96 -120
rect 40 -133 42 -125
rect 70 -133 72 -125
rect 17 -198 19 -194
rect 47 -212 51 -210
rect 59 -212 63 -210
<< ptransistor >>
rect -23 24 -15 26
rect -54 -3 -52 5
rect 57 18 59 26
rect 116 24 124 26
rect -23 8 -15 10
rect 116 8 124 10
rect 54 -69 58 -67
rect 62 -69 66 -67
rect 59 -82 61 -78
rect 40 -113 42 -109
rect 70 -113 72 -109
rect 53 -170 55 -158
rect 17 -182 19 -174
rect 47 -187 51 -185
rect 59 -187 63 -185
<< ndiffusion >>
rect 56 2 57 6
rect 59 2 60 6
rect -21 -14 -17 -13
rect -55 -19 -54 -15
rect -52 -19 -51 -15
rect -21 -17 -17 -16
rect 118 -14 122 -13
rect 118 -17 122 -16
rect -21 -30 -17 -29
rect 118 -30 122 -29
rect -21 -33 -17 -32
rect 118 -33 122 -32
rect 15 -125 16 -121
rect 18 -125 19 -121
rect 93 -124 94 -120
rect 96 -124 97 -120
rect 35 -127 40 -125
rect 39 -131 40 -127
rect 35 -133 40 -131
rect 42 -127 47 -125
rect 42 -131 43 -127
rect 42 -133 47 -131
rect 65 -127 70 -125
rect 69 -131 70 -127
rect 65 -133 70 -131
rect 72 -127 77 -125
rect 72 -131 73 -127
rect 72 -133 77 -131
rect 16 -198 17 -194
rect 19 -198 20 -194
rect 47 -210 51 -209
rect 59 -210 63 -209
rect 47 -213 51 -212
rect 59 -213 63 -212
<< pdiffusion >>
rect -23 27 -21 31
rect -17 27 -15 31
rect -23 26 -15 27
rect -59 3 -54 5
rect -55 -1 -54 3
rect -59 -3 -54 -1
rect -52 3 -47 5
rect -52 -1 -51 3
rect -52 -3 -47 -1
rect -23 23 -15 24
rect -23 19 -21 23
rect -17 19 -15 23
rect -23 11 -21 15
rect -17 11 -15 15
rect -23 10 -15 11
rect 116 27 118 31
rect 122 27 124 31
rect 116 26 124 27
rect 52 24 57 26
rect 56 20 57 24
rect 52 18 57 20
rect 59 24 64 26
rect 59 20 60 24
rect 59 18 64 20
rect 116 23 124 24
rect 116 19 118 23
rect 122 19 124 23
rect 116 11 118 15
rect 122 11 124 15
rect 116 10 124 11
rect -23 7 -15 8
rect -23 3 -21 7
rect -17 3 -15 7
rect 116 7 124 8
rect 116 3 118 7
rect 122 3 124 7
rect 54 -67 58 -66
rect 62 -67 66 -66
rect 54 -70 58 -69
rect 62 -70 66 -69
rect 58 -82 59 -78
rect 61 -82 62 -78
rect 39 -113 40 -109
rect 42 -113 43 -109
rect 69 -113 70 -109
rect 72 -113 73 -109
rect 45 -161 53 -158
rect 45 -165 47 -161
rect 51 -165 53 -161
rect 45 -170 53 -165
rect 55 -161 63 -158
rect 55 -165 57 -161
rect 61 -165 63 -161
rect 55 -170 63 -165
rect 12 -176 17 -174
rect 16 -180 17 -176
rect 12 -182 17 -180
rect 19 -176 24 -174
rect 19 -180 20 -176
rect 19 -182 24 -180
rect 47 -185 51 -184
rect 59 -185 63 -184
rect 47 -188 51 -187
rect 59 -188 63 -187
<< ndcontact >>
rect 52 2 56 6
rect 60 2 64 6
rect -21 -13 -17 -9
rect 118 -13 122 -9
rect -59 -19 -55 -15
rect -51 -19 -47 -15
rect -21 -21 -17 -17
rect 118 -21 122 -17
rect -21 -29 -17 -25
rect 118 -29 122 -25
rect -21 -37 -17 -33
rect 118 -37 122 -33
rect 11 -125 15 -121
rect 19 -125 23 -121
rect 89 -124 93 -120
rect 97 -124 101 -120
rect 35 -131 39 -127
rect 43 -131 47 -127
rect 65 -131 69 -127
rect 73 -131 77 -127
rect 12 -198 16 -194
rect 20 -198 24 -194
rect 47 -209 51 -205
rect 59 -209 63 -205
rect 47 -217 51 -213
rect 59 -217 63 -213
<< pdcontact >>
rect -21 27 -17 31
rect -59 -1 -55 3
rect -51 -1 -47 3
rect -21 19 -17 23
rect -21 11 -17 15
rect 118 27 122 31
rect 52 20 56 24
rect 60 20 64 24
rect 118 19 122 23
rect 118 11 122 15
rect -21 3 -17 7
rect 118 3 122 7
rect 54 -66 58 -62
rect 62 -66 66 -62
rect 54 -74 58 -70
rect 62 -74 66 -70
rect 54 -82 58 -78
rect 62 -82 66 -78
rect 35 -113 39 -109
rect 43 -113 47 -109
rect 65 -113 69 -109
rect 73 -113 77 -109
rect 47 -165 51 -161
rect 57 -165 61 -161
rect 12 -180 16 -176
rect 20 -180 24 -176
rect 47 -184 51 -180
rect 59 -184 63 -180
rect 47 -192 51 -188
rect 59 -192 63 -188
<< psubstratepcontact >>
rect 52 -6 56 -2
rect 60 -6 64 -2
rect -59 -27 -55 -23
rect -51 -27 -47 -23
rect -21 -46 -17 -42
rect -13 -46 -9 -42
rect 118 -46 122 -42
rect 126 -46 130 -42
rect 35 -141 39 -137
rect 43 -141 47 -137
rect 65 -141 69 -137
rect 74 -141 78 -137
rect 12 -206 16 -202
rect 20 -206 24 -202
rect 47 -225 51 -221
rect 59 -225 63 -221
<< nsubstratencontact >>
rect -26 35 -22 39
rect -16 35 -12 39
rect 113 35 117 39
rect 123 35 127 39
rect 52 30 56 34
rect 60 30 64 34
rect -59 9 -55 13
rect -51 9 -47 13
rect 54 -58 58 -54
rect 62 -58 66 -54
rect 34 -105 38 -101
rect 43 -105 47 -101
rect 65 -105 69 -101
rect 73 -105 77 -101
rect 48 -154 52 -150
rect 57 -154 61 -150
rect 12 -170 16 -166
rect 20 -170 24 -166
<< polysilicon >>
rect 41 27 59 29
rect -34 24 -23 26
rect -15 24 -13 26
rect -54 5 -52 7
rect -54 -11 -52 -3
rect -34 -10 -32 24
rect 41 10 43 27
rect 57 26 59 27
rect 114 24 116 26
rect 124 24 133 26
rect -25 8 -23 10
rect -15 8 43 10
rect 57 10 59 18
rect 57 8 116 10
rect 124 8 126 10
rect 57 6 59 8
rect 57 0 59 2
rect -63 -13 -52 -11
rect -63 -48 -61 -13
rect -54 -15 -52 -13
rect -54 -21 -52 -19
rect -34 -30 -32 -14
rect -23 -16 -21 -14
rect -17 -16 12 -14
rect 131 -11 133 24
rect 131 -13 145 -11
rect 82 -16 118 -14
rect 122 -16 124 -14
rect 131 -30 133 -13
rect -34 -32 -21 -30
rect -17 -32 -15 -30
rect 116 -32 118 -30
rect 122 -32 133 -30
rect 143 -48 145 -13
rect -63 -50 145 -48
rect 52 -69 54 -67
rect 58 -69 62 -67
rect 66 -69 68 -67
rect 59 -78 61 -69
rect 59 -84 61 -82
rect 16 -92 96 -90
rect 16 -121 18 -92
rect 40 -97 86 -95
rect 40 -109 42 -97
rect 70 -109 72 -107
rect 40 -125 42 -113
rect 70 -125 72 -113
rect 84 -120 86 -97
rect 94 -120 96 -92
rect 16 -127 18 -125
rect 30 -143 32 -125
rect 94 -126 96 -124
rect 40 -135 42 -133
rect 70 -143 72 -133
rect 30 -145 72 -143
rect 53 -158 55 -156
rect 17 -174 19 -171
rect 53 -172 55 -170
rect 17 -190 19 -182
rect 45 -187 47 -185
rect 51 -187 59 -185
rect 63 -187 66 -185
rect 17 -192 32 -190
rect 17 -194 19 -192
rect 17 -200 19 -198
rect 30 -200 32 -192
rect 42 -212 47 -210
rect 51 -212 53 -210
rect 57 -212 59 -210
rect 63 -212 72 -210
<< polycontact >>
rect -35 -14 -31 -10
rect 12 -17 16 -13
rect 78 -17 82 -13
rect 29 -125 33 -121
rect 83 -124 87 -120
rect 66 -188 70 -184
rect 29 -204 33 -200
rect 38 -213 42 -209
rect 72 -213 76 -209
<< metal1 >>
rect -22 35 -16 39
rect 117 35 123 39
rect -21 31 -17 35
rect 56 30 60 34
rect 60 24 64 30
rect 118 31 122 35
rect -21 15 -17 19
rect -55 9 -51 13
rect 52 11 56 20
rect 118 15 122 19
rect -59 3 -55 9
rect 45 7 56 11
rect -51 -10 -47 -1
rect -21 -4 -17 3
rect -21 -8 4 -4
rect -21 -9 -17 -8
rect -51 -14 -35 -10
rect -51 -15 -47 -14
rect -59 -23 -55 -19
rect -55 -27 -51 -23
rect -21 -25 -17 -21
rect -21 -42 -17 -37
rect -17 -46 -13 -42
rect 0 -78 4 -8
rect 45 -13 49 7
rect 52 6 56 7
rect 60 -2 64 2
rect 56 -6 60 -2
rect 118 -4 122 3
rect 106 -8 122 -4
rect 16 -17 78 -13
rect 58 -58 62 -54
rect 54 -62 58 -58
rect 62 -62 66 -58
rect 54 -78 58 -74
rect 0 -82 54 -78
rect 62 -78 66 -74
rect 106 -78 110 -8
rect 118 -9 122 -8
rect 118 -25 122 -21
rect 118 -42 122 -37
rect 122 -46 126 -42
rect 66 -82 110 -78
rect 0 -121 4 -82
rect 38 -105 43 -101
rect 43 -109 47 -105
rect 69 -105 73 -101
rect 65 -109 69 -105
rect 35 -121 39 -113
rect 0 -125 11 -121
rect 23 -125 29 -121
rect 33 -125 39 -121
rect 0 -209 4 -125
rect 35 -127 39 -125
rect 73 -120 77 -113
rect 106 -120 110 -82
rect 73 -124 83 -120
rect 87 -124 89 -120
rect 101 -124 110 -120
rect 73 -127 77 -124
rect 43 -137 47 -131
rect 39 -141 43 -137
rect 65 -137 69 -131
rect 69 -141 74 -137
rect 52 -154 57 -150
rect 57 -161 61 -154
rect 16 -170 20 -166
rect 20 -176 24 -170
rect 47 -174 51 -165
rect 47 -178 63 -174
rect 47 -180 51 -178
rect 12 -194 16 -180
rect 59 -180 63 -178
rect 20 -202 24 -198
rect 47 -200 51 -192
rect 16 -206 20 -202
rect 33 -204 51 -200
rect 47 -205 51 -204
rect 63 -192 70 -188
rect 59 -205 63 -192
rect 106 -209 110 -124
rect 0 -213 38 -209
rect 76 -213 110 -209
rect 47 -221 51 -217
rect 59 -221 63 -217
rect 51 -225 59 -221
<< labels >>
rlabel metal1 58 32 58 32 1 vdd
rlabel metal1 58 -4 58 -4 1 gnd
rlabel polysilicon 58 9 58 9 1 we
rlabel metal1 53 9 53 9 1 we_bar
rlabel metal1 -53 -25 -53 -25 1 gnd
rlabel metal1 -15 -44 -15 -44 1 gnd
rlabel polysilicon -53 -11 -53 -11 1 din
rlabel metal1 -44 -12 -44 -12 1 din_bar
rlabel metal1 -15 -8 -15 -4 1 bl
rlabel metal1 -53 11 -53 11 1 vdd
rlabel metal1 -19 37 -19 37 1 vdd
rlabel metal1 124 -44 124 -44 1 gnd
rlabel metal1 116 -8 116 -4 1 br
rlabel metal1 120 37 120 37 1 vdd
rlabel metal1 18 -168 18 -168 1 vdd
rlabel metal1 60 -56 60 -56 1 vdd
rlabel polysilicon 60 -68 60 -68 1 pre
rlabel polysilicon 60 -91 60 -91 1 wl
rlabel metal1 39 -103 39 -103 1 vdd
rlabel metal1 71 -103 71 -103 1 vdd
rlabel metal1 41 -139 41 -139 1 gnd
rlabel metal1 73 -139 73 -139 1 gnd
rlabel metal1 55 -152 55 -152 1 vdd
rlabel polysilicon 53 -156 55 -156 1 sen
rlabel metal1 48 -202 48 -202 1 amp_out
rlabel metal1 55 -223 55 -223 1 gnd
rlabel metal1 18 -204 18 -204 1 gnd
rlabel metal1 36 -122 36 -122 1 q
rlabel metal1 76 -121 76 -121 1 qb
rlabel metal1 14 -191 14 -191 1 dout
<< end >>
